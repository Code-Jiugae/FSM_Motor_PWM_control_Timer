`timescale 1ns / 1ps


module mode_select(
        // input[1:0] i_mode,
        // output[5:0] o_value 
    );

    // always @(*) begin
    //      case (i_mode)
    //             2'b00 : o_value = 5'd10;
    //             2'b01 : o_value = 5'd00;
    //             2'b10 : o_value = 5'd10;
    //             2'b11 : o_value = 5'd10;
    //             default : o_value = 5'd0; 
    //     endcase
        
    // end
endmodule
